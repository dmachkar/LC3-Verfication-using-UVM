//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit [15:0] npc_t;
typedef bit [15:0] aluout_t;
typedef bit [15:0] pcout_t;
typedef bit [15:0] memout_t;
typedef bit [2:0] reg_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

